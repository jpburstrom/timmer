BZh91AY&SYY�� '1߀ryg�����0����`>>@�� ��Q@�h � B� �� � 7�յUF�((�k!"���&�4����A�� �44 S��@h  �C@  2dшi����4ɈMi�0����4���4d� �h   *)�S�iOS�Sd�6�����4�4̞�`"HB&�S��F��L�Oҍ���FM �Q�::�*<Y���������PM��/>�t�w�5�8z6�翧կ��ٝw�~?��vj3���n��O3Ø6���HD%�à(�&�*HUI�ρGc2b�:�b˨�J��}pj$���&�1=�<�;q�k�N^�?�ǃ^�熑)JF�h��h
V�*JJZU�
��
B�B�(��(��(Z
ZZ�h
h)���JD�JJh��

J�"�"��#�U# T �P��P� cSϰm�x����,DQ�o��D�̷ٞP� �&���p�l�nٺ5�j7f�B8�UBYu��ml+6Z&��T�R�d�隈CE�����8q�cd�cu�e��Či"^\X�a�^i�B��F���ic^)f%��l�0��8�i��͖��Қ�M`	�,�]dۉvY����dcq]ph�kAfck0m��K�kU���\c,]��h�a�[t���l���7@��sR��L9(C�*P��X���^�Ű[6�e��]1�6��]��e�b�p�!p���l�-�P�m�uр�1:D��M���j�"HC�uVdj����6UT��6oo]k�\,�����x$H�c�K:���4�<'6�,gF/�O?+��[ıU���:��'��Z�9PI	%[3Fk[B,,N����:<�ϥ��� t���{�roDb	�hc��c��DN���ɷsF�J#�X�6(m*�,4�N72�J��V�	1�s�l�m������d6*�t1�E�.m2,�n((V�(&Z&�:Q�����t= P����H�L�h�к5Ѷ��U�75�r�<�?|h����@_p�{��w"bC$N��	���`�y\����L��+M�:3k&�UdT�	(8A��o�2��ޜ^�ܛ�-i*������:����X���۬mj�H&"�D*�����U�'\L�-jNLMH�Fm���df\���EMM��w	]n@�7h��*-�N,��y�"��m���-��o-�6XE-)7��(q-������$�H'V���,NL����N�����k�Yq��$?D\KE3�rQ�Kjե$�ZF��w����l�E 4�Y�IDD�� 
=K�ϫ��mA��x�&�:e����#N�q�{z�R$/���wP0�_^�D�}a�y�'<W��A�}Y i��;Ei� n<��|0�v#����^ζ,�5 ]�$|ڰG��)��}��Fi�<̝�vG��I�&�� �u{uI���$� 0�j؂(���ל��E��$���υ���P�㚗2��T� IL�b@��=dV,�@Ѭ@��@ӤAHEgp=&��3�Y 2 �#���4}��S��Dj��q�����َ�B��=Uȋi\Ďp櫢m>]�V��~7�ْ>�����Xs�ٷ:ɴ0j1�\�K�ń,[[��m�A%��j�Ώ�>���g<'v�)˕�$2���"1&~�_�k�3_Z��46��$Q9����`7;���&{�*�B)b�EKQ*:�bu��"ջU��=c ]�-8��u.VI��A�G/#����%��$8P�#���Z��Ä�B��1b��K!�B�c���xp3bv�*��u���v�t��e��������
X2(�A��/	��F�Ax+}z�0r����@�u{=Iߌ5ҵ����s�0 ���쾙�#"#*#���[ђ�1R�P���aUr$¾�浈��9F����K6ɸ��S�q+b(0�%�A7�V��D+��Vb{+\we]�jvĪ����V��lNDB�;��۵u	�8 �����7���4/��V"v����ٜmU���2�Cq!1�mD����bRwP�b�T�B.�B#|n��WN�L8�0&5C�k�9��޻���_O:����"&Lۆ�*����>J������#+�f����0�i�h�$&�i-]���.bC�f��֓6�vm�e��1�!	��X��4,Ic	���;���z�k,���͘�Ai��R(�M�:��$�uD��{�osE^5�C��="$é17�b+�kobfmd(�D�Ll�@r��f�j���I56�7�:2�U��<ٺ]�Fv9	��>:�zt�����sw�F�Ծ^�l����zkrG)��&��+�+N$r���L8���jr�6x�EnB�`ӫ�3��p�4�vj�Lkߛ�!����o��v�-t�É[��`�Bz���I����F�gN�f�`�LĈw�� Ȯ�2�7*XM�Uhc�8�)lŎܗ(�d"!���H'4S&C)؏M��C諸����������L��#Y$YA%�Y��޼�4Q����W���#�D�&���7$lT>�y�;{{��c�qY�:w"oc;f"��f6x:�����R�ʾq�"��L��;�ZE0�ˮps,�Ȭ�1��\��df��1c,Nc���zO']�x+�'�n�H��uA�]�H$ΈL���j�"����1f-�sU%���Im�ywt龹�E��f��4MY����Oi�}G�����.�cG$^d�����F�l�f<�vv��X:�6�KK�Iek�Uj�a0�m�`��a��]juzIB����gM����$�[ʆ���kq���r�S��~�2-�ֺ��k���j�̪퉪��6l��6��q�����[wCb�F�ML�*�����Z��X�A���l�Uee�&M��z��;����uư��#�2\@�k��J��A*��6㹘�+-N)�Ū"RL�UZ^�fJ�"k�^�nD]we�t�@��蜛gJ�$(��Fm2"PJ����ݙ���F:�Oy��Ff(Y��n4c�W�+	��]ѽ���:�H���M�M��-6�7b�nDGR�f0=�Aپc"+]V�7g�&�$P8�Ԙq	��
s2і��s�3>�	���p2w�u㑴��늕��B'E�֝dS:�8£��:�^��v�y�˙۵pI9�����2'�N
��'eG��!D%	�	�0Wl���Q{Q���F�UQ9�����yaYS3.�jnx��X�B��4-���/���,qtA:}Q<��j˙��dȂ�m��X&�.�Y�λsq�+f�nB;4Z(�+n�ah�.t�D�4[&�e����Q�fBJ��6ͣ�N���Ҕ=����[צG�-�1v>��\�צF���5�u�9b��G�%��N�H`��\�Q<�)�l�n3���*��}��T���n	��	"��܍�!�uL���d���)��.^�S]�8��W��|v�T�5���+��ݕ��3nu�9O6�V�嫙�[X$���)��٠O�ƈn@!0���	'�T3l��U��s'��oOU\�����{U�"�K`/a݅�&��7쫷nڧ9��;ѽXN�Ⱥ����Ũ��	�b�Y���6sD�)�:+��34�kk���h�/2����r��[1.k�lwFkU�Z����uӏ:��!�0Z.j>��3)x���R�ú�n������6+�ǿ>|ɾ �w2�C�ʌa�F��JY����ݷ�47�͜VZ�ekQ��v����t��8�$*HHJ������P�&�㣞�|&�`В�!	�(Р�Ee�Y �� \J��N�\�#@��".PT�)D@d���-JgK���H elE��^���(��)M"� ��Tޥ��U
o����Y�~��F��&�k�x�P  
R����KI�v�g<�����ݳ�+M7�ޮ���b6�$8�g�4$��nyd�tV��a�?;ŵ�1� ����0��ߙ@�H:�B!���
�c�39c�>^�y�'�ހ(�C�� �g��i�| �_�_*���	 Q��#d<����?���q���i;bS��o��h����|(�3�y��=����?{�/6��Y�H�{�'wz�[�~<`a�HHB��9�?�8p����;5鯩����ׯf�M�N^�X�:�(�M%�Lx@�C�L~��_L92���� =R��F݅G�2�@�hX�"�V0�+kZ��yY5ܢ��~_?�^��!�l��U v��$�	8�7��ts��`�V�b���!EA.�9Z�ʋ/�UTzl�u��tC+��^�P�y>�������#�"��������\�a�'X�|N��C�q�0��U��Y�j>�t��0�r��࿓�`s{��R�QUmې��_W�^� � Qv�D!����$�А�l1Y��X�ljJ�]��c������dG=��x^����;X�ˢ�=�Ͷ� =�X3���2�m���9������Fג���)w���P����W��.��nSY����,�4����0�������oA{�|~�jd9y��$c����"���C�6�K�w0�PuP�[��3P��rx7E
��;��D�|?s�o�ýz{�>p��p��I^��C�����G�|F�ƀ}�2'�0��0�.��gN0�T�R�h�$}�>A���@p�f��#����7� {o���w�����N�<��$�1��n]X��@�!2��0���L�.L_G^^���k��0Zu�mǄ+ ��6�\�8�f�j@h"�p7����J���r����2h-"ql��A�UUF�cz/�ƍ�6V~U�fLR�7Ҙ�ø��<��_¼�DB-��ﺓ���;��o����^Cj�������5WWVSn�@�;�ƚ��׸��Ï/Yx�"Ҏ֏W�]\�I9uv��w$S�	 ��i�