BZh91AY&SY~�Q w߀Ryg���w������`�R����M��!$���?2��j�Q�5�Ȟ� h��є��LP�        �&MF&�04ѦF�a!$z�mʞSOB6��ѵ#M 248ɓC�� �� �M4i��H��h������2i�=4��4z�� ƣJ$�m3�I+�ՊĒ�k�[M�	-��RC������wO�l�G5��+����6b ��{�M� \�Q$)�M5FZ�+�� ��!��X�a۫�/+�G�y�^���50;tf��*�/Bw�S�1H�>����u��-ǫSk�+��nFF�1!e(m۲��r��/�g�����`!��dƵҡu�&����`�C����h�vw����x�$_p���cKZ�$���l�"��uΫ�)�=�gꮔ[&i����n�*t�6�7}Nn�8�Jpr��N�U�PQ+�@�M�1���TX�;���b�Y�WP���' ���n��]D��@�7���p�B&H�~E��ˢ�1���XdN�������H-��2vs:��J����U�匨�4UlJ]�, ��%�H�w���ajcKI�Ay��� oΪN�PHI�@�.d�-�B EyI$�b��ЫRr�ij�rѨ��w�"&l4ݬԫж4��cA�65���C%4���ɡ���2C#;��NAT��!�GE��v���ۼ�v�u�i��7m���MD��p�x�D�P��@w���.*.:�A�!1xbˌ�蜁R����ݍ�1E20b�mV�.`�:�8Svb�5px�tM0!(M�H:���C`���^cKTe��+��tǱ�_���P�g�]�����5*��x����WCU
=5���q�Q�$ZE`�W�C���+��Xx�dL�_�UQX�\�>}���ȼ=@�;�u�$mL��	��A ���K^_��E� �"`�A��O��\��O`~�-X$h)*I����v��wX5̊p��E/������f�&ڡ�+`}~A�N�T�9�� ��a�!+|Eٳ��c�e��B����N���ޚҦZb�4��y�SQ�i;Z�JiI�\�
�K�
�C�V��� ��+�-���5&�
�[K�%�"AW��V�Ul�2�{#�@A#\P=�#���A����3��������*I.	bU7�}�(W:��3.���K
���q�[��2ȩ�>Z)�� ױh���%�h�6a�q�8A�40~5�}��1)>���DeK�!�~_���%M��7�_�v�h1gYy�>g(��*��x���H�(:N�^L�+���Oޛ��M��e�H#"<��ʬK�4p8)�I�I/9�/7�9��'�Š��P5|۠�Q���Vbc�T�����|���E#����S2'@zT{ׁ�\�o�:�j�'D
�A"�E��7�,�#^̷� � �9#�D��@� �}�����e� I���`�4�/PmL1�< 1�i%��MXt�X����T�TL�)d`�"����s'L+J�)=ݕ��+�99+˗��Z��,TÉ��q�LB�:�kA�������i�ʃ��̖���@�D��A�Bt�J�,-0Xq�Sd�0�|_�@�����t�ŒZ���W:r^���R�A�2���ʒ��`+T��@�ǢX\fKr�$���M���|#c�=�!��1����]G����H�
 ��J 