BZh91AY&SY�m ',߀ryg�����0����`?�� wp<P= � @( !
  ����Zڒ(�J��"dh�&����OP=MCѩ�h�Phd6�jx�T�P h� ��   dɣ�C414i�20�4�2a����U��  �    �Dԩ����G���ɵ4�0�   D��L
��U?T���O4i&OM&ЏP�M3 jp��Q��EGA���肂hAw�\?/��qF��m�������3�>��<�-�*��7�O�հ3f�Y�@]d4 
0M��ZI%d��EQ���u<�ɕ�[آS�$�2�ыD3�W�WL�@χ�.JT9�BH�h��J��hb����ZP��)ZP�*�)��iiB�(
�����
F����i��J���(�������B$hGŌSA�QBR4	@PR���u�����٧��&��4�eQ���O�H�E����
��7'����S|Fn�mZ���ٳ�&�P�]c-�[ ��͖�I�x� F��Ժ0�f��m"(%f�mDX��X�Cf�n��#H����m�g�r��åqZX׊Y�e),L5w:��`�se�c���Ą�F�mK5�Y6�]�k#q���W\$�ƐA٘��kaR��hn*��cm�7Xj��]5�1[ +����!��Թ�SJ�ʔ :�4�5ׄ�ql���c��Lm͢��b��uز�2�\+e��9�t�2�mt`G9LN��:8g�C� ۛ2LC`�C>b�_7�8�6�Y��yc<�@j���PeW4�3IV���*ڒ�L��y*8���]x`JR��|�I ��gw&�Z�t�$����4�9R��
G��e�rӧ�=�p�tO��JjDa1Ew�=��\ٱHt㳎����tm�A=�	��hg'�c�Q��]��ѹ�Ķd��dijjs2W:�R��6��7+m�-m�)j������R7�Kcɹϛ�u�zF�6�X�f��9yl�"�_�|����?���Ș���vB~�>^W,�}}L˜4��͹��U�SD$���)�d�b�zqzkrn���������:����X���۬mM(	ÄS(�Tw߶J�BD뉁w���Iɉ�ͳ�L�ˑ�^���9���+���]E���Ś�7��//�٩�r�1�v��PA#e�RҐ`�pJMB�B�ۈn���N��u`k*jB��Ȉ���d�B#o׸����C��
�@�&�
�L�$|=�{���\�^"�C,�|$�""P�
=K�ϫ��mA��x�&�:e����#N�q���9D��SAE�$�^��$���e�H#�ב�A�}Y i��;Ei� n<��|0�v#����^ζ,�5 ]�$|ڰG��)��FA��2v��g��'�|���H����'�B> ����b��ۇ^r�c�$x#>r��AB��j\��YPJ�%2�a!r�X�~<�� ���"�@"+~p=&��3�Y 2 �#���4}�!z�uRǳ��c��8o��=F�t*�d�D[J�$s�5]i��
�=���E߁�#�|2�@��)퍛s��C���1�T��[alXBű��)VڴXh�6���9�'sts��ݥ9r�I��D0��__]���k�'M���GN}�ԉ����"���3�!V��H��*Z�Q�u����F���ڨ}g���Ai�S��r�Lb�9y͍�,�A �p�#���Z��Ä�B��1b��K!�B�c���xp3bv�*��u���v�t��e������pTAKE�#����2����[�'zn��1��+��.�^�D���Jח4jۙΨ�X�RJ���g���������!oFJ `�J�Bj;�	�Uȓ
����"�p�EƟ_M,�s&��5��%c�@�$���&��|�ߵ�wu��*=�6V��ʻ\��UTms$�}H؜��Tw۷j��pA�013sA�o	sZh^*87��D�A��8ګ(7e�$8��Bb!ڈ181Ĥ�0��^��](�F��on����qv`Lj���s}۽j�N�}<�ߦ����q3n4�"�Z\�*N�,�����Z�ᦘ��Bi����mM��$1�i^mi3n�� gf�fZ�3���L��\SBĖ0�LA�N��u����.�8�f2�j�B)P�	���sc�c��ew=�7���/�/}�vzDI�Rbnp�Wn������QΉ�ٚ��I���յ�M�$�j2m�n2vted��c�/D'�8EYA� �����y�_.n�T��Z�����[�MnH�5�d�<�rEiĎ^�{�2<�NP&�h��V�uq�t.�&�N�P�u�>C�����)���4��fG%�H$�
֧7"M>�6+:v��0��Bf$C��pEu��I�R�m�C၂&��nK�~2	�@��)�!��b=7�����NVf��s��3c8�d�e��f0#z�L�F+�kw^C� �%Лg��ܑ�P�������f(�܉��혋W5����n+{{!K��*��`�s3���i\�k.��̲7"����V�Ir�B(A(�`�a�����k,����۪�7u�Pc�nR	3�9�<�ڣH�z��LY�n��Ioqv[e^]�:o�pDd(ٮ�VqG$��S�sR�^���E�h�̗���m�Ǖn�ܸ�YF։ir�,�`;j�U,&m��2�1�'��N�i(P��\��2��$�[ʆ���kq��WNU�y;o�fB�Z�Y �mt���IfUv��v�6DbJ���MuѝE�t6.��od��Ȑ����-�0���Ŋd��[`���(p�,�2m������;���/gq�&xH�r̃W)F����6PJ�����f)��S�eqj���7�V���������׷�]�q]5�:�:'&�ҪI
 ���[L����4fDEYy�T����(R���;��F9�xⰙ�������[�U`��&�얛
͛�P7"#�h3� ��1���y؛��v(h�L8��J9�h�Kx�9̙�t�q��;�:���NDu�J�Ρ��kN�)�\��Q�O�d/��;n�<�e��ڸ$���Tcř�'m��㓁������"��x��+�sz਽��dg�`˥���pL`[��32�v����t(�CB�[j���-�br�&��'�z�Ys5:VdȂ�m��X&�.�Y�λsq�+f�nB;4Z(�+n�ah�.t�D�4[&�e��9�y��^�s2U�9�m�b�)C�����s�`[b&�}��\�Ι�����G,U���d���I�IT˕j'��9����y�8�^[b���J�a�#��`�0!a$U;��d>���L�6�%<aE��Jk��]ת��ώӪ��^^%r�����r�mζ�Nmj���W3���I7�vS�S��@�	���Bad$�I���3��is������W.a��q��wH�����wJޓ�A��U۷	�S������ެ'Md]C��v�b�C�I���1	A�,�ta�9�{ʝ���g5�����w4	ᗙ[�\�Q�H�s[b-���5�6;�5��v{j��ǝVp��5.���Κt�sy���_��m�O�3<]}݊���ϟ2o�@!̿��w�ĬҖf,e�wm���|sg��)Ah��7�!�si���7$��c@���Gg���]6�����^e�ܭ�˒�,�&��gV�bbT�
�$F�P� P��)wD���X^��DR���E��L`#�hP���W�3E�AD0�PP���=��J��)/0� ��j����-��@$ �P$�@��&ыJع9e(���]��0����W���
R]�Lr_TP�����j�z��\)G�9fv4%���O|�aJ��&�D��U��DH;�6fT9�_l�\{e��Y��}aBa�ʀ(�Q��3˓���o�����"=k�`����!HX;��sjy���f�H���i9D,��zk��8U�u/@�B ���x۸����?EقS�{��z�N��]��y�@x0�d��s�{�Z�ܰI+�v���!V���E��/arx�`��p�4��b5�npH��Ó,��^�
 ��@�T@�.��- 7	3$:ɤ�rd1�
I��0^������9�d�� Z�L�$�XA&��'�k8��!��8�3g�
J���V��6�|��)P�1��=�P��=/��j>OAތ�����˩4�Pu�w��P��rM&�:G'�8�u��"K��(�G���A:a_ѵ2��kE��I�0�c٘mK�p"%��<7�w^r�]�� �5����R�����r��a����t�����-��Tm�
�n(���x��������q���QȖ��u�\WFT$�H�8K���9fd�U|Y��Qr��)��MP���B�u���r��X3؄�af��H�����.2�zBUrp��U��pL��q �&x���Y�"�KhA���蓧F�>~�P�s��3(x���q"������������:���ǐ|�������]����8�/Q��d{�H�����D��.,t�,�B�%���F� kT�$Xx$G� �Xs��:n
!�gv+���7��>ë����ǡNQ�N���Kdf.|�����0a"�Z������L�W���j��:&�ġcp��c"�jJ�A�j%�IX�ᴜ�΀(�EP�m5�	TS�-�w��H\���86s�y��[���׊1�3F�M�@c����Ms��D|��g��|}����oX�/�M$�³H,��׵d^���eNUBm��$_2�f�G�X����X��vg�|����и}�@Nӂ�����)�8[h