BZh91AY&SY��D�  ߀Rxg����������`��|���x8< a�� H
 PfA�U ��2 M)�=4OQ�       d)*z&@     �2h�14�@��`�M4 a�H��i��Ѡ      �I���JlMCOHi� h *H����jbO��j<�@�4&G�q芫HAԢ+�y�(�� L�H���Y!$��%�3�����ُ��ã� vy �uD�B�3���9
�4B�J]Psqׇ��9�=M���c|���ї�]>���>X>>1����GN�s�8���	�u�/:�ܼ���u�65���4vx��V6q��:�^�l�����[yq��;�y�ާ
�\a�B����^�:�w�mUv�<8ɝ��Cr�M#,
W�e��6k��:>�!��$��c��׺|�h�#̪�8�IϝXC�ET]$�#���5�Ln�З㗢s��Q1��Sٽ����w��c��.�o_1�
��R���BR�Ҕ@��@�)AB�4!BR4�)@��HP,� �_��|ڑ,T��!������'���=�L����:��;toBl8����n�p� ��t���%$��B'�d�RW�1���2�HA�LK�,�W���ͥr˶�m��g��˶�m
��'�y���k$��ۃ�H�6�hF��ػCg6��]v����ݤ��#lrBM
�s��oY��ڻv�m��B=��)4�m�Β������b��w��_p~�=����[��� ��LOa���j
	1̐�(l�w>�7N��ko5}�#sK�VZ1��6��2@+-Y-�DHu����vGS��>�O<8�5ӟ����T�U8`j�d�w��qkS�E$�3M��s%Ke�$�I�=����雡��PP6ni��&X�-4E�푶�F��O������3Q^���ѓ����v�o���+��q�`1L&5�XOkp`cr��4f���.6��w�^K�+�`k����n�6�Q�hK�����&�����gdv��ß�Bؔ>/md8�����������d� �*���X�
�Hw��c0�S�O���Xhs �}6�S_�	|��<����LO�/S�Ja
�D�N� ��fK�m��rӡbS��"�c��!^�����5}�`龆�s� ���I�Ff$"�j���8��.�﷔st5���'i!@��tN!̤v����ןT���t!�d	�@�1+K_PI�'C�$��l>#���Lb'�R%^fCOBa�%�B:C�k��@I��oG�4�#�gadQGHj�	�/DAa�qkبg#1a�To�r
�J�iZ����ɣ�6��槢 ����0r�M�
��I������]Ir=�b�6� Ն.�[W9���v42��cN�V(�G*�"�d��g���<q��%�:�y�[��7$����ͤvYZ���:M�]�������O!���2����~P��U��8}+\��_�&bf���-�g�l@9pdޝ�HV�D��ȥ=(L�T��<1�p��VE���6��p�U��_";A5(����2`�.�*uGOdۈ#�MVE?�{S^!�D��LZs�uOz�P**+j��&�&xaA���!`���(� �K3vW>=f>��3�6gX�B&$8Jb�$�jr�D�Q�rpfE=\���f$a�ܼ�P�����X�_U*�3��ku�{�9��d�缢6"��9I<:D$���R�� �5�b{0�ּ�A@B�@xY�����0��u�g�sw���`�|�4BRS���n$�G&�e	��W ޓ<k$wZY�OB���ꐷ:읆-�_O<�����_��,�Ή��KL�ǀ <��r�/L&=���>�3�}�J��qr�|rB�\��yd��M��!}7[ڧ6.����6Գ_�_�w��y~��zǙ�O���,�Z!��BD;,��n�u�l���VʂQ�����O��&�n��3ÞD�4�0���@Ǣ�+�/��� +4���w�(.T5����x0��~�T�;�*�e�Y���=�FøfSO�oJ��ft!�P��μ�3`���f���ݿ�43���tס��p�<�#$(�
cŀh���˧Ó��W��PA�x#8�Ŵ�k�k�$�Л��GL�(������ ��ꒆ�bD���3ʾ��"j,ד��Řh=0�_�s+�(8��>K�fs�o���j''�33wp�X�V�Ċ-�ú���)fiB&�^��<�@��-���*���ݐ 	O;�B��i�TT��KF_��Үy�b���ӈu	A�;?�멞�Tܹ'PH��X<�W��s7}z�ۘaQF�dN225$$i��rd;	fv`+$	���-9q�����|�e�lͳ�D�� � ��q���]5�7�g����]��F�]{?����,�����Kכ�{	�9>��}���	�y 	Fp�؈x�y�:���Y�;o*xt��|<���&|�S�0���H3�����{�"�ܐ��`�v���d�Ll�n�u��]4e���WF4ɵ�ǈ�$�{<��	z$�(��b>���z'�h�c�"�����T���;��*��Vz��m��M$'�$:���c:�~3e�#��H�ژ�K"8���Ir�^�Ur���]n�v��A@�͞�S3�s^�1���
�v���������*!(	��e�s \lȑ؍�Z� ڬ�:z��zw�^����m�m;�Ԩ�[[�oj.�^7֯����y��qbs"*|/q�K9D:rC��q��^���pT�j�˚"��95Qv1#�5gC��o:�J2hv�($a�Y��ue�Ց�s�)�H9G��̟�آ{j %���;�2�M����9ä<� �9�`��US؄�@W"0x<`��xa��Cۇ��(p�\_.�U磆&�B��tĒ�̀���
��v�D��6��1��2�A�$�`���B!F	0fo�5d�bE`���&H�&�s2rd�f
e�b�p�4e)���`3.�>8w��*]���2�����tX�
T�J�UU����n���գ��[���پ��(����>m�9��=dG���G�\N�K�-���k�r7����f�wpk��/ze1zZ�RIu�3�+�~��0S�g�l�=�*�hn��Qc��W <K�j�8�>��ꓝ�1��AKGr���N��7.ާJ$vu(g�;UQx%𙀓��c��}<�Mʅ������9I�L���l%�Eݫ�=��Yg�a�b���mm\�F�z�Z\�������`��x�c�~�~�1izV�ד��y�I5"v��3��(� S�m��Iv��Qjx��*��3��֨��vÄ�Cd�-RD�V�����:�Q����{�C�r*��i��9z�o�UM,e���T�G�	��y�x���O��h:t��)-$�&����j�>Bl�V��.�K�˃&?YM��^5h���c>޲�i��S�����M��Jk���]|����rIkl:�)P��g�W�Q����Qe�oc�?��{�T�&Z�noFy�Q|]gh),�e|��4�F��0��~�XC�C�4C��9����d�95XX½}z��prGUyÃ��Q��
�Q#����_7DH��b���v�q0�p&�$�%���ˉT�w�k��+�k�{uI$Io[�pw��RO%�.5vO{7���K��I��k���`7�u��y΃��<9ʨw��5�#J����*n�&lk�=�5T]MrcRwq�;�Xw|�!�R�X<�#���:�Qp��b2)����|�D�f���4�f1T���{�q�nr�RMak���n���oq����y�d��f�
��f1�.l�����ٰ��o)���[-����$�%���ZʱM��m6�L�&���6�ʫ��i4I;�����~�c�c�l�0��ݥũv����۲����V�kl>�i�'ߧ����{�u%=3�g��iq���no���:�{Dc/-�݁�.��?Tbѝ<�w&�	J��T�)(�)'QÌ6�w$S�	~�KP