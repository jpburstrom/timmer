BZh91AY&SY\C �_�Py��g߰����  P�:�Q�B����&�	�i�4i� � 	)��jM6� i�  @  � ��(ѣ�����   dɓ��&	�F�!�H����4КBi���M@����4��H|(A�
�� ��ρ �e&�D0����7 yM$X4"�ط��5&
��=\a�y���A-��9���*�ˤ�Q���91C��҃o�$�6��ܸTfB๪E�`���u�5+��W�
�D4+�HC��� V���X���P���n��.����+�#V��S>
�r��X�,HT���d9A�DmEQ���-*���_��j��������!fѶ���5zL�L�W�p�;I�$�~�-zI�bY���!		,$�I D1�a���Yr�B�H�m���hZ��9r�RTC-gGY�@��c�v�R�h��k���i�cYb-y���%^�%u�cJ�tˠ��N0D�
�AA��H/N��aY!�2A���%Z����AR��^65t#��^���Z��� :VS���
A֝	"H� 0Ծc7����p��<[eʑ���R,�4�h�v�*��J��芰/��{nr�(%��w1�1��%uDI���(EL!�#��ʁ��b�1���N%��׀�}�
�I�h��ꦪ��Y5�TO��H�g�:`ҌHG1%����^f<1��(�!`c�u��G �m(�-#*6�i�V�����3���������ñ0�ŀ�#/�:�4X=���icE��aFI��@��hd�I2�V�����]󙠘*&N�D	�/B���xT���-!h�сX�*J@��X�ӝ}GI0[�����~���=����Fu [��f/;x��H@���_Ȭ���ԑ̘�n�A�G�W�
����U�"�+(�\6Jqh $�z��*����6���|+\�MB�9,�)����fȍ�!H�����R��G�ә*J����R��~��Z���%z�kP�Ku�������U+a�<4��6��E#VQ�g���)����