BZh91AY&SY���� x_�Ryg���w������`޽��6��u�NMt�v�a$���=��*xj�Q�6Q�����2��<�A�J2D�Mh�� 42d��bh�#0�0MdhjD"z�=M6���44@  4R�I���`���� �  ���������SI�Cď(  ��+ST��ǌ����̀5�^��D�!������;��6h�����թ�K�S���&�B0�p�n����Hq�j�_d
��<X�^�V,wj�˱ۣ�l��H�ja���fӪT3�\��5'�b��==��E3�NAv��Z�l�\��J^^E��
ݹ{�aZ���SeU�����KS::2s��un��ѹ_=��L�ޞ�u��.-��L��<�ˡ@�ï2ih&9	�>Ecz�R�U�=�ig�tY&Ĉ�z���Y�I�2!��klCh��XV�Zf꤄ta F���&}W�vI�^ܓ��qq'/.EU���*��b*'U��c�U�][�� ��r�S2G��A$���w�]��Bɢ�4�0��{7į*EC<���k�8\��KJF<TX��C��%am�u��xKm�ł�$f�"DS��͸��o�ӱ�8�1T�b���ʎōu�4���+>�Fa�m�U`0k�Z�-��|\{mP�ky�[{v�Uw�u�|�[y�p=�Hl���Ƅ��UTꥷ�f{xt�OjCD���E�Wm.��};N�ss#LcԘ�5k5���X�UC�UY،�!$py��1�(�d�d&��% ��"h���	1JJ�Q�U�RW����褤b�)���)�%D¥�);�Z�ev&��JE�2�e;�C`���^cN���,+���c��.�|`>� ���-��+[lJU�����%U���
=4�氃ԣPI|��u^e�A��m?Y�ͳ"���ʪ�s0��c~��M���1!��K,>�i�C�^˵-y~S�-�����a<�j�5A��P����'i~^wn�׍C��F�D��
�	�^�1I6ԏ�����d~e/H��s/�B�ۆBW��E۳�s*�	b�t�K��F�q��]�;K%�n!��_:#�FS���d*��mhBւ}T*�X4}���{@j����w׎GI�B��iiȺ�B�*�y���P�����k��Q@�g��M&T>X�𼫼9Z�����,@�Y�+�9y¹ԟ2ߐ�(�����n�=�l�B����`.<�`�4g�h�6a�i�8A�40~u�|w��Ĳ�E��������?��f扳EM�����]�Y�\v���e���Q�L�eĤIj�8^V�ն�i��&Ƥd��@k�ST@Y(yN�ʂVj�*�4�[F�UBOIA� ���A�7 �+�rdK���҂+`�N$�XT�X��] �X�wA	޾r)�B��9]�X���ݳX�@���p WB	(.�ɽx-73�7X��dj���H���l5ʣ1+�ĀB�j��2� K=!i{�A�0�N@��Ʈ�Y%5���"NNAN�hZ�� �3'�Μ�+5�)��[�"�!Q�����wݫA�`��P96���.T���?�\���([M�V�C�2t4��Kl7)�AծrWx��`r�M���e�v%�D:	��u�-v����e�М�����)[a�2����r��_)S�b@���XZfK��FVX����Q�E�������Q�]�2��ܑN$=��>�