BZh91AY&SYD!�~ ;߀Rxg����������`�>]�� � 
 H�c#fP��$�i6��OJ��覚?JS'���h�T�@*J��@ @   2dшbi���4�&&�h �Oi��Q�        RMOEO��h�z���h�z�!��0�$���ҞMe=�L� �h����-���FòJ�Q�T]Y���T~-ՊU�����3��?x��%�OU�����$���h"�2����o�8(�`8�џ
�iHwŨx8�އ�ON������=][u�k�$�� DD*� ����^
ꝳ���ؙ6�cߜ�p���>ګ�������TfAq3�Q[�0���f���M��[6Zd������8�n�
ivõ�m!���8cGd�v�+���DMb����Am�k)1ƢKn�j��F��2��ԡw0��ƂJ��t�<�q���%��.(�4ƻV� 1Yyf9����
�������i�4be��[ujL�Vr�P)�����-����V�x!!F���9y@k��ܐ 0��[^&^���o�n��X�f HL2d�	:Rܝm-*8�H�����}KIU*Zc����եXF�-�f��.غB����;<^�r����g^��ى~6(x�� ���|ʫCbP�69�G߹����u�WB��Qd̒���IB�"�̤�U�	��Q����P� ��Ɂͪ���4$�ȉ���ݿ"(`�<^������*^����C;ϲG��� `�Աg��hiTI���ȳ䚉b��	Y��_V4ڏ4�#��<�0�!%H@>D
�i���AP*Pa�(��y'N�% 8����Du�"J��$	5�H�C� 2H2�Z�f�� �Xr����)��Z
���:�i�b3�P_G&�
$�Y��~V $�Z�[ڇ�-I�P��s� �	7�_�(�B�-�S�%�ea��m��Ch,Ýe� Z␀�dC��c�c-�&"��{w{Y�s�{,�r��ݜ�^�F�FOt�X��٫+�^	ј�3���P�.�-Qy�l8��WUn�S@�
��{[RgA\:�D邖���=�F���T ��a�Ȝ,���3�kH�7%�#fEtힺ������}�f��Z�#����5a��J�aep�\fZ�ޥc�,�Չ�Ku�E��Z�9��Z�=
�Cwu͈�.(��A�Z���So��u�]1� �
��itt�mei����/6��:�Mn��@���aB�١���Z�s,��l����`J!�F+�@D��7xq����{^�݌������9��2���USG-N���Xd�;�/�Ն��ד������=��8�]n�z�뇀�n�F�)��Y���M�dK������\ؙ��\yp��vY�}3ܳ��5��eT��W��d!#�X�&�yF XT��W519;Р����q%�Ȍ��>��
�~T�W��73�bh^�Y��pH6�Y�ڭ���C
!4��M^�]2���<ֻCf�dt9�� >���Kfu�]Y�l@~>��m$�B!6J:�nt�ZCQ�6jJ�6�����BD��-���#�Z�t���P���Osz����ǵ>bĥ6��@��/G1�S!C�T���k���7�uz��^8�L�jS��ͪh��x����l��*�S�Q��W1$(��ʨ�vӋ��R��̊�k±B$�5��ҥl�x��U]Cj�FR�w8Ӊ���4�x+��Tv�QkD=�f�0�e �ī/[`΍�3)�挧ܒI
���or�EQ3y�"��-/e���K�u���<��)q6�A���μ��:t�N�m����3�[^�%ҿ$��h�ج�����W=�F��<�oЍXG�4D%6�!ەSN/1͸�p�_�n�+[w{R&c���]�l�u��BH��17{R��yp�ua1"� -�b��t��|#]u9�Kfq#}ov���C\(m�V���pu,��«�ޔ3������׈�Ve��Xݙ����!⫩�U�F��>���z�y���*z�#I�|�1�e���ݎSk�a��{##�2T�I�4��bQϸDG�����{)��E��!�y�/A�X���(�����@n�P)P�� �E@�P ����L)�Z�n�	�lpԳ�D­`�!m�*H� (�#�:_m[Ei��ן-�lx/�r�`h�_��?~�íI~��z�-6��w2�߼�?�xfk���L���z��x���*7�$���>����GGA�����"��S�!`�����O��nN*!.pB�����f�(x�P�(�I���~������-�Jv�/ض��9��B(�-�w�b؍P�q]�+�';�("��E��m	�����J��=���ӴF%ń�8 81�y���D+���
�L0��xu�}��P4$�wA����Yy�uOo+�F-G����L���D*N15
y�8��Q��t��!fD�p� �.��,�
k�O<��9���кk^]I��^	�H��0j�D׺�1��!�Q��b@�W���9uy�B������vO4qD��%����|@0�!N�v�t�c�)�w�&����7̄lB�j+��A@X�Rw�[`n3L�2�%��UD���o�:��.�U�X��dŸ��&Q#(2��@�è懛��YɣXwlQ��0<���`:B#�B��g�u��`����p�\A`8un�hm#�wq�>g�w����s��s���kG�p�RАa��6�}���Hu����bl:6��NpЃ��)W�c�t��vW��'M�E��)�
k�8���``W�.�71t/B�H�QX?�SN����0��;@�1���-��IH ���A��TYر�8ݘ�n+
�p1�q1K.�d-��끴����� ������b��Z�F�%�n�7�pȞp����ݯ����"�A�I�.�K�"�H�
�?/�