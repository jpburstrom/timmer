BZh91AY&SY�sc
 �_�Py��g߰����P9�A  -��	���dɓ#	�i�F& �(�dSĠ       ����OI�2i��H�  h9�14L�2da0M4����$�MLS"fL�Sj�D�'��l���z�W�W�H��I�H����G��K_��W'Ҙ*����I��T_j�I����IH2T>��2�ҡ۪v�m�la����ǀ3e���2��[��4�������ݒ��6�1q���CQ����R94Sǩ[yoɚbSC��S�ڬ�T�V�Vqq���n�[�4�X��#tqS[��e6_"M�kUg\���}�߶���(�%J�)�o��S�����7�ԳWAJ��aR�3�;>Y���Ņ��s�`a�TTT��Qm��_����R��8e�:�a�I��cU���4R�eJ�PqޕB/�	Z7��Qo����ӒɈBo.�r0�+8��[!�|�
�V�,�ŰԺ�&�6�����m��J����j
D�O.T���U���衆˅���Ju���N�jB*��Ȕ��hA�V�\�RO�/#au����K(eS��^eH�J�ңe��[~�3���[�wW;i9A�}���|�U��<�@0�pc8t{�8|�"�%����>���<�Ŝr��,G����Ǵv�4}m��yeD�e�Y=q�z*��8p%��R��p���$���D��0>�:�����UF�Rӕ�Ibz�Z�!}IT��.qd.�Yg�e�E	{�$�k��ݴ,SA\�f��X�Q3S�L,Љ�$ˊ&�[�\Yq�f��KS�}Q����U.�v�'GT���o'ZM�0�#g)U7`ۜ�%��2_�����`��(�,�a�j�rzRuc�}$�ҙb��/3���NVwrt48˞���*pmr�����3�S�&��TW����y��p��L���%��iơ1>�b}�*
�t��O5JG>��7LRh�Dq]�M�0KӝIK,�tJM��J�
Y/���N2�0���KJ��W�P�"�`���)k�&)-j6���c���̊�pI���ӹ����L�,�_w��������l.#�7��t��q�y�zӊ��K���J����%/���*Pv{�ybqO]���SVoC�	�sn�2SXH�5u�%��)=��p� \h7����E`�Q	�4rr�2)�PF1,�\��j�99�Fҥ���uo9��Mٙ���%��E��ס��?�,�\��O�d��f�s��s�?���H�r�eC3��,TS�c���%!��3���H�
nla@