BZh91AY&SY�Z� �_�Py��g߰����  P��` ���2b10d�2 h�00	H�jL�CCj4�     )�H��  Ѡ@    q�&LF& L�&@F �"A4� �i�$�'��4mM�DH�Ą�(��K�1 _y�$L���#�!���N �i"�m���q�0V4\���9s�h�	m��8 �D�k��)�ME��'�D�t3�����8Ä�ae
�H�Z�_t���yC3)����f�f�d��B)[�M Y��!�z�>��o[-�Ɔ�[;�I�í6~[!���+
@�f�N�t��,q�	@pu��T�7�UEwK0�{��<֌U(%(9^�&�
��M,VCLXAlU�+����\Exѽ��0��(��UT$�`3�܊D����x"�eI�sDC<���&�Jȴ���2��H*ȁ�x2H���	������3��i�sW�dy{����ٞ��9���S�3�����t�3�b2	l��3������
Cjd����%�j�M���Q\`/�ˍ|��v��	{ЬA��� D�^r���H7�BH�;�8�γX#�<��?��l��TA��b������C卋���w�p��mEp3�a<�=%"EZ�ڟ�&�'8J�	(h0�&^ȫ%"$x�@?��q��~*��(r�T׀�i2�&�s�����Cfj��Ȱ�Q�B�ۂ`ҋ�F�Kt��+<�u�� �L�@Q�ǀ�ҤzICYu#��E��,Ր��-1�g��������_��ĘK9������:�1^3i�t5��Z��7r�\Q��Iq9�--�d�I31+Ƅ@`�	�t��D��H����L�,SEYІT�*�C/�iT�nE�OV=�;�{M����-n�s{Τj�=�S9��@ih[� �o���WLMOjH�&4�H8Q�$w`���2Zv-i�aE�ʊ�D��@V')�C�ٲ.B.
���4 jˢұ	�$��!-,���
�T<�$��ɂ�Ơ��P$��AqE��~���"'A�[Q�j��^0��yK�jT�����L�I X�A+�����]��BC�k(D