BZh91AY&SY��K] Y߀ryg����������`2����   .x  ����h-�F 1Z�l)�3Uh�J�m@�H�JkTi�k�42�#MY  C8�T  �  ( �<��Q)=5@  �C44�S�)D�* M42hdd�� �0�b �L�F!S���%JHhi�4� d4� ё�4��$�	��24��=2�M���ڌ�oHM F�J&PɁ0ѓF& 4o�:L�E��SGj� �?�"7 (kPA[�o�>EC��^ (4��Z����獰��~_.3�pW�Pp�~��{ݛ�M(�E`BHBA�D��P" �t�R�T�b�z ��u�ňn��+�r!R)�9UiD�=����$P*>ݝ�<k����9r�y'o����tl�K���~�E9�B	(��TEJTD@TB�!J����R�*�(�UUD
��� ������*�AQ�Uj�ڲ�	UkV��f���/7I�)���v˽��V#��40��\�T�/������<�9��ʬ��+99Xr+�pʪ�0�aFg9��"
�#r�"# �9AYUQXVr(���9QȪ��ʊ�#�VdQG"#8�QQTV�#
�dG9Y�g2+��(��*03��FfTG"�"�8r�fp0��9��xEx\���G�����o9��׼ �0��"���\Ȋ���FUg+ʌ+�29�APAÅ9'+#g3�AY��9ʣ��3��s�Vu�6�ʈ�Ps�VA\��sDs��#*3���eUdG��3���QU�G9�VEg0�eFaUÙ����"*�"����A�p9����ȮTdAA�&�Es2��̈�s��FaXE��a\3�Ñ�8Ur���FW �W3��29U���2���F�r�U�9����Ȯg
"$��6�xDx��FA]�?NyÞ_5��?ϒN{�9$p���ӯO�^KaIxlL��W��K(��ͯ��rw�A���xE|~����fs6pv
����sX��鹖D��"W]��ci9]t��������P0�e�a�*�Vn,i���,W1sxƖ��F[It�eea��b�,%�[-B����$�Yl����f*�t��2�يB�Y�[���:fm6���X�f6�Pl6Y��T��lҔ�	�6�ڻ�h	f�&%�9�Բ���-[�L�fY�Q�#ct�f�靆�pr��!4�bD9�-�������.��K�la0�]�n5�� dҎn�`ՌԺQ؄&-�̢E)�j�V۽V����x�̢��P�㩿.�{���l3Ms����ӆ@�kS���g-�x�~o�{��uN{�Ҫ�"���*�u�""D��'�Sz5�g;9�d���i����|��e(C�j�f� �Yt�/��S[�6���8��Y���si�L[�@1���(a�ℷ�����9����w�ɩ�v��.��k�0��b,�Xm��Sj�4�d�c5ڙtm�c��ȐΙZ�6-��n�-yk)��5䜜��$�y����)�	��I���{e�,�Ù�2c�Ӛv���	�1af��?�	}<I��#�:nL0�J�!7ą�:�t"����0�����A�?&Q��N_V&�IY�WD�0�(�K(�br�
Ɯ8P2���JBF�C3�#Fr�.�YV��CL�jH��!��3���=w�m<�����\�D4	�Tؘڒ�;+�sS�L��E�u�ه;�A��ݥΌ�L;���1D\��W9ʚ�B��,�N8��ѳL(;�"䥥P�p�I�bRa#,��W�R�L��-2�����m#�Ɩ���<�V~zz�%ǅ�Dt��&a����{O1���xP�B2�4�\W�3�6(&1nm�OS���,���8s0��ȱH�)#���P[ͦ����$�{"\V"�1*!�]\�e��Z�m�i�m�9$�7�2��0��A�I?�"9�W%�/u��޼X���Ww7%�#׋+�~����_nL�Ţ�:��"���*0�w�0�Tp�:"���6�q3$8MKS��*ׄ����
� �*�����aQ�+��~�ۼ��]J3YJ�x5���,1�---��--4.�-�aj��U�^!e�s$[���#��:��ke��X�����i�DeUR*Ҟ"��,>G^�+(�YZ��Q^�%����Y��8�4"+--��eB�&XU��VQ�eO*С0���zs[Q#X���KqF�:��oV{��)P���ؖ��<���^!�=��r^|��e��e��#HS?�#p\g:r�I@X���7p��ZkI�m�Ҋ�ܙ�����y$�:�Į=[֖�F�K�a��A�=C(i��Jߝ�b���*iE9(�+h����Ez����Wq\~�|��P��F�cH�S�Z�y<�̹E�.�
>,E`�<P��I�nJ��*H��/��S��.$��r�x����V��K�z�-a�m�YiűԷ]!m�2���+�u���O��^�J�(K�[aq�6�[�A�u� �1�UeX��a*�A���A��#��XvY;[)^ٍkt�͞�,3qb��l��؆Ƒ3�PZ]+��x���	�L�a����]�x�8Y����[bv����(���(��1��~)~?W�TY�,��Ŗ.��H+����ض�J�Z�I-�9���"ťåx�@�����d���E�X�$��&P�<a��x��%���0Ѥ���	4��9��d�z�f;	1I,љ�rD@�4�(��R3��$�W+ύt�D�P�!m�&�!�B��(D��\4��@x:A�-�i���$$���3��
bTL����:["�u�M��-?#N�$�>[ǳԋ��Ku��^��+:����6�S��u��G^8q�t�o[q�7�)x>@�.ie\�F��a�6��4�3Yq8��2��P�%y��BSn�P�I���n6P����$�Zb�h�i������=,��ęi�|�������n���t�hI{�Z�U�RR!%$���m��q����*�ng�.&:"ԼI��BF��4~��M?dh�,��%q�r,�I	cJ�	|Yфx��$��{��a��
<��Fe�#J���a�Ȟ��g��c\�k�+h�H�k0��m�]�	�y��I����g�0���cm1t\�a%y+(��t��:`P�,�E��	&�.����B4�E3p��� �a��~��%)�SQA� D�\g���|s���g���te�͵�ZIfrJ;gʹ�",��IQ�����ݓ�9��ϔ��;.�a�Sk�v�DF�Wj	��#]���3%����֖e��O���ٻ�x�,uM�IDB�,����*6������F))<A$�7���"�y.�i��I�J�-B�� ������#��� �rH�;'H$�Q���]`J]�J\�$D�%ړ��R1�Y'N�7�l�
d���ώp�	4�tTt����s���0�m�=|n}�!-Z],�b��R���	���l�핥��E\A,�6R�պV0�m5���<������!ֆ����n�͘�t!F]���-�Lar�3�2�-�ml�k(P�L�F]ky��4���c�j͈E�m�I�,ҙ`�+R�l!x��>1���L�,��l��4��e�;������xH�f�\����<R�mP>((�H,�*1���Z~�S)ӥ���ʣm��������>i���fb%"�`�a�I:��|���S��,�$�$�8�֞0��6�F||i�M4�9�s�Fm��_&\I1%%�#��5�C)���V�v] 38~���p�a�N�Y�0�?��}lC�#��!�����8r�m�f%�FQg�8~BV#�t�(\�-i�!-<Gh�:r� ����4��m�b��2S��J ���s��(��4��/%�_I)��ܻ��2����S��ZL8��K�p �\XQ�A�(�v�2�D9)1MMb�BC�]�a3�*�틓K����q�׬��ч�id�t��>�����p��(�>�E��dZ�I""H\��uh�˖����d�0��n0���r�J��S�-�[�3���`� ���NI*����w��u�֬���瞖�-��_i�a!�� 6vQ�ByѺ��P_���(���40��jZ"�,��p^/��_=����g�@8Uef喖���2��4����IF��4ӎ�4�q���8�ӥ4�DBD�)Ƒ��ZGC�[g����O�Mz/�_z!��O��>,��M&ؒ�J	<Q�I��t�OZVI&U��/7�јD������s�aiR�sĔl�#(��]0�]�_T
"bP`�Zt@�i��A"7q6æ�Y��| ��;(��?2&Zd�Ը(�n�#�l�����+5��ɔ�èH���#�I(�]�ݖ>�Ν�.�RL��*�>9��ÆYki���=�4�{�^��&11.	0�ώ���ka�����a�.A���J!�ˉP�C3E�Y�a�m<2�7$��U�>���b%�%IR�Ҥ�u$�[uǼ󶜗r�c��z�ܜx���il:�.x�v6�	�����n��9���[`�q �m�\��iV�4�D��d��EUv�ԇ���^��k\��2�"�e�B��A�Vf�U%lVmu��*6��#m�L^|��K[b�q1��a^K�aj�Ax&6�p�dj��E����� GK/���$Z$Y�J<t�R4��{�Ĺw�%��4F�0�ZE���-
Ԭ����,���`�G�3��X��3L0�Eٯ53:a��������M��R:�ƛB���p,,��0^�{����0�Di⏹��|޸N5�d%��3"^bk4Mej�e�ZT�U�D
��Dݤ㈲��s��Q>�[o��$�:i�$�o#��/��(�_0��](er!4��i�>i���$����a�.L��ն�|"�K�
���e1�Q<��O��J�I�3C��GL='�QF�|adx��I��ԼIF�d.�}�V�Q�f��3]+�3BS3	$�����)$�p\����,��=�[I�?4���+�dC;,�D(�$�j��i Z��F��I��w�Ό�ԩ4�?���<#BϘ�Q?;�)Aޮ$Q��<���%մ���B0f`Y�I&O����z� ���	�g�σI � �ΟBXQ�o8(�,�^�R_t� c��4	�&
Qș"e�p&M6�ϼ�0��I$�ȶ}*C�e�֚zÌ>�}XA񼒊���%|����R����6�=��mT�F�8ˬ���s�Iv��ߏ-<|�h��ɶ�����3%$$-4�N��h�I�((�e�Z]0$��mi���l��m�j�W)���[�e�,9����4�Ü�D2L4��n�7��PCp��w�t�O�E3��n�UYӦa�g�>�B�|KJN��}�֜,f|�L/�'�u�����{)U�%EI""D�H����d�/~�$'-Sd�du��$�xPi�4�(Cݮ�QVh���[���L�oZw��>/��،����6��Z���Q�i��f�c��3ŝ�4W��q�O!/�	g������cIr��fr� m�P[���\M��Qm�5y� �3���xo�]�Rv���Z5k��n�!B�*���1+Y�2�%D%�6~K>�$çI?@�s�z�c(��0�)1��
0��(��$i�O�$y)<x��wó|3���J"<m��m=�����l6�M0��%y(0�y�$�9�z��,�I:`|�bLгxp�書p5�����e4�%$ͥ]CQL@�	� �4�I}=M�E
�I"�c��i/c]ie"N�Xʿy�E�i �/g9�KHΉ5�<#lPQ|�$��0��O�#d���,�Q�t�U3z+�RY���$8�$��y�E�A$$sƌ��,�	Ҙ�%����̱f�WVZFX�[�Xka�0҄a�KŘ1� �M(�u�|]�ꩥSn/2E.Wh�������%�%D��.$74oQ�x�k�\�a��DÆ8GK��袺�:h�aܷ3�ʻհ�b=�w%S	[�E=uIͮ��i;�66.��b�x��v�DOr�1��iMb��6S&�d2�k�e�i�|���w/�Kf^��,܈�nj��ts�.��v;�\��5Td�m�]�ս���qm%=����jn-:�U��Eو�Ml�8$J�S	]��Ű�so�v]�Z]��wqz_k�S؜���=��3��1f޹�Z����/j�}J=o���{v�!<��Q(¦fKԫ3�v�Um��+��M��u]�Z��n^P�q��3���{'o�������ú��N뻣23�Z5曳�;-ޭޗ7mT�Ԅ��Ȃ*�K�jSˈ��LR����H��j�M���8�{՝2b��[���;�eʈf��]P��r�aӣ+EC=�U��Q���0�H$d0�9f�AΘQў���x��s$�� � ��t�1���6�Y���WJV���j�3�`�4�s�!��ԕ%}�D4���t/��s1"�}ҏt�x��$�6�I��i�p4��&`����	G!�g�	�s��(���/��<t���vx���㶖"�g�:s��N��^��s*W:���ѷ�T�m�]:��L<d�B�k,���0��Ia�K,�Ώ�
�DC��Y��,���Oy/�/��!��N�i�Đzңq"BH:&t(}��m���i�t�Ǎ0�t�pk���=����H\*Zʘ�_��i]�6����GT��0��ag�~�!�v�}�BH�TD��2I!"x0)QlJ<�B��+��ԥ�\O/�.�W'��ve��L��"`E5�h\\HP��0�Q�;[<8ȅ�A�`�؀�P$+1J�AY����Y�yx�µ�j�DR �T� d��Z��d@���.1�J��(�j��C�m��EV�t�h"��U ��
@X��R�P0ƌ�i�ns�fQ�C�J�]cպ%�JAad�AA�2���ղVߍ}�c�g��^:�+_�(�)u��tU�S�?dn+���>xIy�C�����7W��U��h�)�Q�>�p�wM�����4-T!�N5�ZUY:3��bu��얼��kw�[�k����7$��D�t��<�\���F���d?�'z��c�^)��AaR����98�V����% Xm���!�w�f�h�90��@��xm���7����_��@6^�Ā�:�� �2�ܷ����T�y$�-M@t��S����� �p����`2�n�*3:(:MAp�]T�$3�����T�N۬��?���a	�����  ��1椰�����@f�2���*�t�b(0���Q��E'���pC�b�V��ƀ���拟
� >zw�dZX���6'�U v�1d�B�8�Ys���16M�d:<�C��|,�Q�>��L�7�`q��D���t�cl2h� �Բ�i���A�}g|�H{?�=W����qpt��,�*�.�t��/7A���P��o��R�˄�a�Q�>ކ.ĝ��}���ZBI7B��U���we�W���38b���t�0�PP��r���c�i}�a���.˰İ|D6y̔�<]�*�K*�N@DA�C�p$S;�~��I�)
�4��v��O{�[��@,`��]�*(>X p��U~�l�em)�1.vR*��x�)M�髞)r^�ZU`�&�L�K�ȧ�K�޷��Iu�R�����m{��8��G���#A>���5ͬ��1Yի�����̠ס������^�BAO]_d�s�Q?���oٻ�9�~�?����c��K�<�]4��r9�7���	j}��aH��'1��96��R��<�"���~��8p�/���$D�ܷ�;��/Mģ�~f�g����py���y���6ᒜ���*�q�.�������`KK���F�)�%�|"\��Nr	��L)�Ӈ� �4��K��d[���+�������Ȩ�3DH����m��J�/[�@� �7���P�����|�{v��p[A7�Ld�ϲQFe�W�;���HV��-�L}+�g�AN��(����Q��i���Ҧ�@4I�׀`oK��A���(����������63� ���J|�F����㻸�k�ZQ�wy
^�	񄀾��Co�rE8P���K]