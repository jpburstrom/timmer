/annex/objects/SHA256E-s4908--8dd73743c8acbb8e980c1d806faefc4dc25e0051426436f9f426195bd3225f79.sv
