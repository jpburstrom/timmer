BZh91AY&SY�1�f J_�Py��g߰����P~�jT��4h[�A�ɓ&F�L�LSSS�d�I��z���j�@ ����Hi�=O"4��A�=@���&L�20�&�db``D�	�F�F�z �M�a4z��LOS�bX�UPZ��/��%�TRi���\`6!oBh���Ѹ�R�Y!� 7��a�0���8�4U����v�kWc:��C�\��{@+9��0�1%9�#r�P�&<;���9���}LJ���&�&8�U�5F�2=&��i�2M���9�cE���,Qu�_���|����ތ0�Dr�j�R�N<�i��uuaҳ.�UTu݅HmY�C#��ZXP���1ʆB	L�M�]	��di�(d��{bH�j:ҧӆlq,�[Bl�Il��ɳ�T�^m1i()�/��34K^��A��٢��WN���W��x��p��61�,m��i(C�#gh��f:J�0�`#����㉸�q>$D���v#$"�����P�G����2��f*�8��R
X��4>���cY6T)qh槚��+�[֣AN@M�s����t����$�u��~�g��������3��y�d��fT06�����?�|e{T�|�#��#ҚH�bl���J�������-8;�����H*0Z2�v,���9�i66�Q�1^FBC�X%�Da�q�
qh�,SDJ�s3#�2�nClZ�BĆX"e��5TB��x�O�)�i|D���@ъk-8v7��Q�w�� �p71U5^��qgYڧENl�VLIy�;�Q�����Au����[��f�:�&�C�(a�Q�y$�R��50�
@���H#�Xy������A$SK� H����$!����G��M(d�H2�r��T,6�A$��H�6A#c念6�j��e�"~�"�YDb��C��4`�3������xplݨϤ�*/��l5��	�� �q��I�(/3�d� ��{<�t�d�H��Ά��`���!�9��Ȏc�a�>�S�b^v�
�C�-Y+��3o
��Z��'�k5͂�ѫV�f��+�5nd���1x�ͯ�R"MƓP���|��%����Q\P-B@��㖤?ᓘ�&��3C&�Si����b�nkt��9�;
#���q���w$S�	C6`