BZh91AY&SY��Z� �߀Ryg���w������`�^S�0��j`Y P�Di6��=%?S��cSb�<�dz�4!�6��5=&$�P��     2hb14`��@	��24	����g�zL&	�S=щ�bhhmA�L��M`&i�L� �DH�4dL��LiO)���#M @X���q$�?&(B
	$+��@;�ܯBKb��	��m�o}�a���L��?W�8i�{@�%��#Z�\n,�� �bi+Ma�������F�,�4ka���~%ɧ~�hB=,#������S����WŪ����S6m� ��Q������nFF�QR�N�FS*9L>](��gB��x���b  "��tKggM���EU�S�oT�'Aǖ���)P��%=!5XǕ@I �bJ%pHA$`8�uR|���Z�ڥ�-]X�#x�1��Lu�"���T��h�r�9����X����&��j���Р}�'��7eK7-u���|����F� pX���,@M���2�-�v߽B��H�u�඼[8��6\�*\��Q�v�m��A�F/�{�|8�����%��D��C�]B���Apbf,�NZ�-(z�ͪ��*%�*���%exf�`��8�d#��t�[8ciQ�R�"�P2�P�&�)��T$�BM0�$,�+BbD�F%��4�3��*��0yY�2X�Fv,�jRa�P3\�1�!a���]���'xo��1ʛL� �q��m��I
��� ��f�X��͔�w�Cvb7�Gi�EgF��l��>/F�RF�1d�L�1p,��F鑒��V�4�md��E�64`�D�4j�A�75\��!�160���'<h�ǆj��,;�׉��u�?����ϑ��������ϑ�V^:�����Fpr_p�e��z��m?9���Y1m�B�Ra+�މsJ�tf]��3��uJGE0B�M��(8���j���W�\5��C 7�H�pʕ�9C�^T��Vq$�w����6�`'G�a=yJ$<~�1D�I��g)Z#��d!�/P!�^>���PgF3�*M���K3�8���22�S]�
x�[x2�wV�V�U���<��j<$��M"!�/k����v�f�u�}z|M��.p���`H9�wW�G.)���ai��H�� ��ޯ�����\SU�3�<h�A(�����u��~>���mXH5B�XiR���g�o".�ͼ�\jOy�o����E@6z6ʿ�jeQU�>k=���k�Y�yq��yY�Zi���6&��kON��.$�^_�CY�|�����*�p�q�_�w$43�Zy���0-V1�*�����e�P��yݐ�]m���&ƨe�@䌽�@���AC�:�*$��U�_-�NBH1~D0k4^W�:hj�b�����r�Ĵ�-f�y}q6J���Bw�\ً�3 �t��U�m<5�V�V_
Ǿ�f	���
V�ɼa�-Wo=��k�zE�`���;�Mi3��E��@!L�n8�:$��3ΈC��5��
HPg}��\K�V������8#24��h���CS2tk�T�`�Vk4S�ҵ�Ey£F�����v|����,K@�ds�aS �R���t��q�.w-f�E����NFB�@�ba��!���4����X,Hۡ��j�.��(#'A2��yx���#X�k��P�aB9?�Z���փ�\cX �`L͓#�zb|,�nQ	�y�X�v�^q� ��{dJ����`G����H�
��U�