BZh91AY&SYZ~� r_�Rxg���w������`�Q� �k�
V���@5�y*�Ju�PD5)�S#S�7��5=1#@Sji���j��@T���� &�4  ��*��4�@   ��&�R�@��     ��db0�`!�M0�!�F��D��Bz�M�O&����Q� ��CN((�äDG3�B�L�,b//[��,f�,�\s�}�?���˚�;�iZ����Ơj�����Q�E.�^)3�P�qj.�:�l������_�]�'�XC�!"�H�����]�)�	�*=O2����H���/�v0m�=<Mf6����� `�.���,��4�[���n.3)`A��YE��v۸��In�k�lP�U���łP
䂲�0͚�)mv&��lP�1x��.�q�f���5c�Q�2�n�<xـ0�a�)JcMu�������-�v���8�L#y[R3��ܮC��t�ƕ��QSN�����R}+�	$�K�i�	h[~va�r��U�.8.M*�B� ��00�_p�{�P�������x�ŹԧJ[�`5(�P-�����4�`C��i�z�ݧI
RwS�QI�uZW�-���߿K�V��K�.�!��E^P�.ڄ0�9c�~Ohz�w��LEk� �!qQv�aʃV�V��2t�ޗldx�lVi��bwLa���LA8�8B�]��������S7������	 V����.��J�r��j���R��]�vDa�B�J��U$���,r��3k���ĴG6�����j�B�<�l]�䥳�JH�q�t�L��O4ry�Hh)^Q��L�mG34n�(�K���VE�_MpF�
R�nEгODsN4(��� "���+�| �8@ͣN��>=CX����6l�īoR��K�:��m74�Q����b�K5n��)˦�����t5,���"��g�xi�ܘMc]���2�|(E:�%Ը��Y~ΐ�^�ص�s�ڈu�-&;���c'�4A@�P-)�[:ޡm񳕽;*�f'y��]����鳓�5ğ��H�23�$�񎢪k�sj/3�](u�",x�̍���-�O�--��+�'����
Gv�D��t��d�����Uq`ƭd�@��H4U��ٚ[��D�oTV80�T�.a�e��ꫩp;�F�f��
SKE��%N��˼�2#*s�)�Є��T�����%"7G�w2���mz�Ѹ��]�ס�J+3��g਎�w��HVs��Q�Rު�xӞ͡��ؐ��Exy�w~lP��|&�f�#b+d�*�z$�y������ٍ<�X������)�з��f��\�GEq<w�.�>��/:��S�ȴP2����J��N�"Ӎ
�uMIvH2�ol���I�e�z�	
�N���.Vh���I�͉:�s*��kn6)�wL�!LO	��+�D7k����]#,��IQ��H2L6�F�p���5i%�,u"B�liY���jU��''��wp�V��C�̂mn�M�^!Ww����س��;'��`t8�{z�ʗ�V�QYnהּ�b�3�v�܇5�o4*�o �f�舆RI��s��w:�/���9�pIٍ�rawuVR���_ޣSȅ�&fk�f�\rԔ�o;��z)���k����H�S����ٕk�b�se#����x�2��I3w1]Z��S졺+xٔ���Naq��գ�q9�����]��p"LA6)0���m��y�L�g[��l��w�IJ�i(Լ�s9�{�^���|2�oD�h��x���ڳZ]|�����HPD�I�ݩ��A�w�EF��U1��Em�I=�����e�;�v�e�!���=���|�M]�.'\m�/cfl�p�x<���0X�l�;/5D*�lt��H�z���v����{W;S�G�gfK����2�|K"����g�ciK��r�.z/)̮��W�W]<�]v$1���N�.[��9�4��.c��='!!�D$�$��(Fģ��U���|q�Rv�YI��bK�!4�Fz�Z��EG8"6�:��DfKX��Q�"QT�+r3�PQ�M6��wGP{6ټ��*uka�-�H���"Hm�!���i�W�f\�T��{jå<��ȷ��z7u<<�y7�����\Ud�]��ש�ū��f�9T�j'y#����+1��'&���b<���n��|r������N2��2!K`����O]��~�����2�4��1���C��R�O�C��3�9��n�kgy�L/yK�wm�c-�Z��vw��&*���z��U9��:U��.}.M`�^�[k��-�M�"`�H��+�	R�Qz"�s@2�cd��k<7�@�y�c#��\`y���t��<44�^grcM�E�BK�Y�}z��P4��P�K�j��%t�+Jz}��wH�R�����v(Ak�o�k=��G�/%�T'���F\���f���>��$G���X,���}��4W�f&hA{�q���'V��3
,V��k�v�sa��KrR�� ��g��&��3^!h�Xo
#�6b�PA`^˶H��F3��Fı^���ͱF����>[�yu0&��]��%��H�]��Yj�!��$CB�T�K]���%,�
�0(���f���ļb;����H}���rf��_ؾ��oe���ٵj�����9��qA���:���ҽAs t��O��pU�p�
bx`_�1��c�80�}!��H��-��<�}�]:�G9׃CG��5���GM�տ���˸��T�`��MwR�ن�DV(�X~9̭QBdL	l�ӓ<�a��S\��Ѝ7��YI��!iS�ج����E��jz�$8(�F��aX-�s�/߭8�H�f
����K_����p�
��Tț6@*� ř/��%:�n�o~Xo[H9�dE���`[̸a���"�(H-?Ѐ