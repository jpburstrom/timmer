BZh91AY&SY��5� _�Rxg���w������`^k���s-w5YWv�D"hɤ�I�0Bzi�i���6�dh��j)��#@� 4 � ᦙ�&�`L#��i���!M6�H� dz�P   ���db0�`!�M0�!�F��H��И�&M~Sj�Q�S��( � �z�� �L�$����!%4	A�����Am�O�Ɗ����n���ev�ʚ]X�ff�MF�- �7n�F��Y5w�x��p]��in1bѡ��>�}i��_M_��榛h
_0��|�K�L�7���Os�lP��R0!�w>ܵ�Z�bSp�rpZ�1�V��7���"�H���tE�7���1%x� �'ځT���M����-;/�U��bT�6�U����$�1��pG<���A��lmjz"e�TE�)��	S�����s/���{�Zg�I�����6o7��1f��N0F���I.47/�p��r+sk-Ƽ�慎S#j��˄��MU���v��b�`�,�YE�V�@��V0��xj�����T�%�������)�h��╢$1s-�ZQ�X0���>J������6���p����cq��gd@8t6Z���k�%�)�|wT���8�%U����LX��1�!�)���҄�·v�*�(w0�Ձ�a��H�EeLYd�J ���]|�߼l�x��uw�\r(���=-�Ow��T�t����4�ޚ�keGFG�N��r���XH�o��wJ�����LK��K#}�+k��=<A�>ĸ���4���&�I(��WA�?�w#]�&#�9.�����v���n�T���������u���m{����F�D ����m�)��Uyi�"Xx�N�#
�M�QT]|\x�\�������m,rf�\���%���刐U����[C��U+������.�A��	d��d)F�����t&sh*^k-(� ���ϗqt�7���t��L)�%��X����~t6�W����J��@��J�v`���	t�����O��f�1R�m7M	��h�Kj:�c�:�7l��� 4-i����{������eBDƗ|hk��ka<���I.=����Y^ƺ���y�2,G|�+�̩%�^���i��M�P�R�T L538J��笚E c��]��6��.%p�1N�Z!�s�<�F(�B$`�hi�T(H�73¨Om�RԒX���(A����4͘�f��<zu��zVL���(�ڙt6s8d74Fe�\�[ r$��g�i�����ID2̲1��CC8Ӄ?�1�ZIҀDc��j9��,,Y�=ar����TJJ#~�n1X�(���k< IMݓ���$�-��A�B�b�Q�X���9��I1��u�Y���Ek������$�e������ۡ�r󬫁@�V�Q�K{1P,V�]�&]}	��Dr�W�ӽ�K/�X�-�A�cb6XL�逬�m���U���������!�`c�0-D���rE8P���5�