BZh91AY&SY��F8 _�Rxg����������`�|� �z ʂ�� H 	� ;ށ�M�F�	MA��iOMM4ji�P4�  i��z�@i��J24�0�1��q�&�CL	��14�@JaDSE= ��d     T�)�SG�Sz)��d� Ɛ   �"&��d�z�CF��i����h4��i������z�����@��"�7��ش��oh�����<���r��s����z�WK�6�}��"�G`��Տ˥KC֘�K�	8��"��Z&�J�
�m�l��b���9a�PإR4ӂ4%�F��D�����ﾐ��1U�,89hۈH�*oA7jC�������(qD�B�z"ǚA�p��R+y��l�L��j�4:���L����B+%I�"��V����V5�o�	U朾�xǕ�ܔy 
�'�:�8���� +���duCl��������q�1�uM�=�޶n|��2���o����2��)B�-R�-4� P-"�!JPP�-P��!JP-!�`$XbX7��x��igJpo^Z.N�?�zl�vs���LE�qH'�֤�"�#TMQI"eJ%$�TblN�(J;(�n֩X�qR�8���$뱴K`�"7G,dm8����k��-�[kmڭ�'-��Y�<V5Q@�-��eq��u��l���br�Z�S�([,��Y]b���-mثi!6��&:�+$�&���YlR[+���+c&*�5pu�m��V�-�M�i>��t�𷫂��)K{EBk�L��(�qS5嚙KL���Y������ө�|\sj���$����Q��K���g�f` ܝÐI�f`�����sy��;!ġ��8uu�P�R�t$�r���W�:�TQRH�4�l�I�*[�PD�A'�"�Uu˩��PP6\�	4�R�CADQK���sF���v�'H�,�L�Wg=�9�X3=Ft�]���k;��t�,��7B�L�Z+;��i%�	�Q\μ��0���m)��D[X��*hvZ"�)j�R�SMH%&�u� H��6��\�0����"h����d��`U��7��+�!޻��_'�JS�M�	ǳ e�_Hp�!/�oI�w��Q��?^�=5B�Q:�Hgl�2n[j6\��������I
�^�`̄�i��M�5FS�BwE'89��E,�n3� "qe�]��DQ�����V5X�4C6Ba8� ":�@O^|R{}Ї�� �1�K_)���t:rK�P�C����G��%����'�9 ZS>fq��0��!!ݵ�_ $�췣�H˳���(��5K�rSFh| D����Z�*��X{��[�V�p�p�A�$�=^��X��֧� ��3��k���~ U!I2мY��R\�D��;	�a�����kb8�]9΂ �,�gXІ���(1���<�$*��j+VD�M�6��R ���n��B ���D���m��6����<7D+��U�E{<S���|Ƒ����v���1��ږ����X�{�)�x1UqJzP�����*��< b�,f�a�P�tB�z�Ȏ�MJ&o�`�#&%§Tt�M��C������-��C��!:����Sކ�8��5�5fs�3\9_@聈bBՏFC\ -�� ̚��n����#��n�3�}	ӈ���$�����!8�Iu\AF���S��~O�bF��κ�	�M��ń_T��3��ku���~�P�M�{�#^��9I<:D$���g �7vk��{0�ּ�A@B����� �1�E��� �nb��/Uࡌ�vE2(��8���d�q֛�2[�uڜM�Vꥍ�,�tp�L��^a���p;���/�����7E��'�#"����  ����]t@^1�缹�a��c��V���P\�Ǉ!!(�n��Qw�3Co��"Ϧ볅�l��Bm�g?T� �%�f�DK�̗���'@�8<(F!�n>Slh(ˮ�e�d��T�<'���$���68�"g��H�T��Tk�Ƞcγ��"����`d�I;�A�*�GTW��t��(E��R0��ۆX��|C�{ꍇ��V����ںbxB'�,/�y�f��o��EYk�hf����C�
#��4x/T4FHQǋ �uC	�O�&3����]B�**jZI�E���J�h����P��
�:^J� <��+�# �k������'0�y��� *�n�WNe�Pw�v�a�-�MD��fn�K��y��Dr��:xJY�P����*�?��-���*���ݐ 	�6�,�-3����a)h��U�3�_�9zq�! �3�z�g���,N����4�x?�;�Ⱥ�	�p@D�dI$&(�B,�	�S�2��K3�Y M<��iˏ�=�{��/�,ͳ�D�фD^N7�9��2*���42�=[��`�6���f���^L�d�y�1g��s��|�`����	�z 3�GDC���9�7`�Ω�yS���]���)��!w�ϞjxF �2ay6���\�@=��E�iT�ꨒ�Tj417+��	+���cI�WZ#��k)���X-W����n16�j��-�#��j��j�D<�Ax0�#���D|��sv���V{	����������Z�lY��y�f�/�G͘�}����#�� ��K�v�⫗ߏu��ڎ�6z��纯_�ڎy�uZn6v�F�kü���'O�n,�o�"DlOb6Aj�{U�gOP�����Hb� �H�-?�`xLL�Y���	x�Z�SW��С�3U��x�wg(�NK:Y��"t:���pT�j���*lpr2hT]�H�MY�P� ��ιҥP4��PH����U��VGtu�bFrNQ�|0y��݊'��BV��
dZʳ�b��ɳ�8C�3H$��%�
�UO�	� �������3�xֆc��@��k;np2gV�v`XP?�6�R&%)$'�i���X��{�`� ԃD0B�L����׌�́ka$V	Y��d�Ri�ɆH�`�K ,��a�L�4� �����*|Ԛ
��.�aeZ�W���ĐR�%JU"����}�oYK7�^�H|���������i���ɾ.}���h���z�>ީ���4}�/��U��,�fw7�lnѤ��]�����x���5�G���.����rG���Ɲ�c�{�s��%?�)%���?6����_O$�a�`'����I���F��49�&����)�܆s�	'8�s	>4��^���К�T-;�xxY��bS/�d�ʡEݩ���$}�@�����ĘC�֩&�me�f�Կ�L,�z-�<�-��ũ�Z��^LJBE�I<�#)H^��Ij@^e�uU"�K5�*�S�������|slT}���ꚢe��E %D�p�~}�Σ�p����Y͑����|˞a�#"�h�I4]'1;�j��60^9����^2��A��Z�%�$�b�\�mW���cգ�y=.�6,>r��sT.�g�'��ƞ�!SJts��c0zt*f�$�͑�������o:I��9JR�ExN2����E�-�����l�v�Cj��y�I�O��*�^*�ގ�d�=&��é�~v502�u{c:(�Ñ��Y������*�4�y'~_V�r�4I8B��+�.�^&L�a��јk@��+���;�F��!�f�b��`�082�	%������v�<ϣ�Wf�(�	%z�C{�ꔩ'��.5�g���}��܌����;e�Y����^�t:��<��T;�{c�!N9����.�C�=@��8I���2�g[�o�U'/J�S�ZJ=ݩw8{c�KI<qϹ�K��;��P�gRi0��*��d�/w8��YjI�V��rg97�&��J��8��ɺ�sU0��s],�ɢjd��2�?6m�ɧv�I,�m¥�)�v��ɓD�]Ue���Ꙛ�O66]�ֳbo�n7<����4��85��ؼ��Ҙ��ױm���lI�?ק9*r��]nD�O�{����N?u����v�yثM���@��LΓ7�,�G�l5sh3ld,�%"�J>B�r:�Co�rE8P���F8