BZh91AY&SY�`s ߀Rxg����������`�|u �9�  ���� H �z���� �� ��	��Sҟ�LO$ڟ�h4�2P=A�4�T��L& F� i�`�&M�&�L�bi�� ��P��H�426�2F@h4 B� ��?&�� ��   T���d��M4��5D����@��4�N���wAEw�@��h70'�i!$���.����x�M�Ӗ�`�S`;Oz&�y͡�}���L��r/|�]QQT�{�U��D	8��E�J�5�֮�gc�BU�,5��8�F�pF�i�#�!�H��۳u��qx��3�\�Ó��BF��G�R(�>���\�4J�)��,y�5����T�޸���	$ɜ���&�T��e�XF�h�!���"��V���f�5�o�IU�?H}#�l'��N �T�O��L-Uc#�I1�;YPك�� n�ی�/�;��i����j����6����wk����7��ΠR�R��!HR�Ҕ@��@�)AB�4!BR4�)@��%��	a�`�sמ1v�Agzrq��.OG����\G���N�V#lؤ��+H�H�TRH�R�I%��
��$ۃu�V2�T��B&��	:�m�1����N+er4Z�q�kV��v�c��kv�Ec��TE$KclY\m$��m8[-�k�������-��WX�c�K[v*�HM��Ɏ�J�+I�c�V[���J�Ɋ��F�q�m�A��KmuZ;�����\!U��+6X��L��Ae�C�� [1��FH���+�p�|7�8�I�f����M��[���@5_6LVߒHv���]������vè�����<�UT*T��������:�-�:�TQRH�4�6-��J���I$v��
f]�͹�]$	+��ń{⥢��"�� �f웷!c!����N����3Q\t���كI�g�@�6E"��H#1)"��K��:"�VzQ��-`�)�x̟�ŗ�P�f�#v�਋k�� �M�DV�-V�V�i����|q�$ٙ53�ˀSL:��F>:�'�8i�?�X~�M�|
�Hw��c0�S�N��XhW0 7��M~(%�M�<��J8~'�K���T�'BwI �풦M�mF�ː��bS��"�c��!^�����5}�`龆��pHN���3h����p`N,���;���R(�;�?� �	`ia��	`�	��t���@Y=y�H	��B,#�8ƭ,u|0��{	���/C<Bh[a�h���$����d�>r2@�����OBa�%�B6C�k��@I��oG�4�#�g9,,�(��R��њ700��بg#1a�Ts�nAZ!É�iZ����IzS,w���Uő'���Z@I���R�-Ő1+	u%��K��L���V���O�z��kN�;�u�#!X���1Pc����S���m�ڊ�U�&�bM�:Ԉ#���ӖHD\(�Z�`�����w��n�<�qD+��U�E|}����Q�t������_�D�@���v��6z���9��mԤ2%��U�)�Bfڦ�qU����@̺����m�"���#�R����3ɂ�p��=�n"�ফ"�<��o/�N�A&-9ف:���q/Tkx�N��\��w@�1!�FB6 � �2hc�m��ǧ̎��glα�"�LH�L�N�r�D�Q�nl\짫����Č;ۗ�u*ܛ]{���S"gwD���o��ޡ웼��F�Q�r�xt�I�(.)����n��e��a��y*����+z�1:bF���������0X~vE2(��8���d�q֛�2[�uڜM�Vꥍ�,�tp�L�凌�4���!�f_=Uy�|n�5�O�FE-3�< �7#Ⱥ耼c��ys��\-`��9��]7b��<9�	�7m���������g�u���6rЎΡ6Գ��_�wފ�3sX�%��K��U�]��B#�)�4e�Y��E[*	F�ӂm?�x�A��3��$l�~L*5���<�:��/��� !6L���Ar��ptuEx�L/b�_�U#�L��e�QY��9����~���oُAe�_TW�D�T"��%��8�l�o���Yk�hf����C�
#��4x/T4FHQǋ �uC	�O�&3N��Ȳ��\�5-$�v�"��ۥc�TQhu�UG[/E p y��V1"FA���_]�5s^Na��� T~�̮��,�w�v�a�-�MD��fn�Hc�X/7(�VևO	K3J7��E@���Ԓ`�X��T7� H���e�i�TT��KF_��Үy�b���ӈu	A�8x���3��{�'PH��X<�W��Nd]{�e8 "Y2$�<Mclm<$Kp�nd�:��y�ӗJ{*�Ɇ_*$Y�g���9�,�*��o�sNdUI�heNX�#ܯ�/ͦ�����Xv�ד5�/^n�Y�'\��_,�'i;�Bx�� ����0��y�����v�T�=:n�vp�
f{H]��3皞�5��^M�u�7Px�m2�T��Q%���hbnWKrWE�Ɠ���G�R(!b�(��o���<�gl�a�����1��ʑ �d �_�{�">Hs��SY�l�=���َ��B}�tHu-w�,�u��3e�#��M����Y��C�%�;zqU��ǂ����GX����=n����W��e�G<�B�:�7;[#s5����TBP���7@�ّ"6'� �tA��Y�t�̬�OL4�(�1$�K A"���������ʍ������55}�`-
��5^׀�wvr�t䳥��2'C��\NI��W1$T���dШ��ܚ�����7�s�J�i۠���gg�Ֆ�VGtu�aS�r���̜Ԥ���{ƣ�W�|%��V�o�yMЦ:�b�����VɃ��"SL�'3#,�ܮ���"0䝄i�P�%SX@�m�R�bԄ���l���&1,�� ԃD0B�L�����~��3 Z�E��Vdb �"�cI0�����2�90�&iC,�1V�Oe&EUʗb�����{	�'�e$ f(J�K�l�Z�Sy��V]^Z�9�^*��|:܇����a�R�t��QG
l1�0*�����4܌)T�-�8�A�{��`�Dz �Xrp����ԭ�x����;>_�����������.����.!��̜l8����w)1`:���L�s�M|�䧏r}�h$�b�� $�����>og[$�P��P�z,��1)��[Ȣ�k�?_꥖|Xh�dœ��ع�YF�f���KL��y�<s0q�~���R��19�2�����*�Pha��F�ƌ !ɤFc�w��1��Ie���$�<'Xv;��	��@J(�V�5�ZǝG(��Z���3���+��704N��UM3�M�j�2=xL`�q͗��<d��NG,9N��KI���\�mW�y5ǧ.ó�9�X���m�gD.�m�'��Ɯ�
�''Nlf��S��ժ>��|z�z�@�jk���Q^��+Á���s8��1ѧ�j�s���F-���d$��$�>g�T��!ʗ�i���>�WZ�1�<�����M^FTa��t �`��h
��G���m��tr��y!�C<d�&L�a��0��](�m3�am?Q�4�A,&i�uIe).u�*��ﯨ+�[�h	%z�G�s�䔩'��.:|��:��ڻ���v��c���0�N�خG!�<�����|>�Ԥ������M��с����D�1L$ɕ�2T�jηy�̪M�^�P����{���a��I-$��fSoskGi��Mg@�m�КLSII�K�V+q�Z�d�B�6��ͳ��KW'V���S^�QA��5R���N�k�`m)��`���l�K-Z�e�l]�a���f�d]UR��z���i�e$��˲:VjMݛ�ŋֻSM���-Kɽ�])�kJ��Kk=��RM�>\d�}�'�u�5=��yW����|,mn���8F�Q���wvx�[��1�-)�����=V.'t���B��Hu���H�
,c�