BZh91AY&SYL��� �߀Rxg���w������`޾_5�24  �׵�B��	$&��F�4iOMM��Ȇ4��hdڃ �?
��@4h     4��a4�C �a&&CL� ��
TѤhd �44 d h"�S�zG�i�4h4 �z�   �2�d	��	�C@ G�ɏj,�D0h Y<�d�a* �T ��-��I$Q���~1�ó��ڠ��=�3�64���j�/F��R@�$�QVk�w=m(`b�f���㢝Nf���M@9&�H=����=Oy��[b���е̐��Y��R8��u4吲!�X�nXۑ����Q�!r�N�P��XbօemЪ��i6�,)n"��F��C�B!1�GKrIE���wYBv5������(ݧ�uʻ��7N�*1�)���s��&8(-h�G��T\����Ⰽ䖪I	��h4�!*�G��_��u�*N��E2׷�$ cMs�E6�J���d����5���Pr��b��V�\vJ�v�3�x|��B1�Ɗ��g�B"Oo�^��O��7�a"�j��'��!��݊a����Wn $k&�;US4[+5V:�,�8H��{�5�@w�F��Q�g�*�l�#��m�0O!e�u�a��WF�zFME�X�X���0��X���Ze�� ؇mB�~�k��[[{���Ո��&�ֱ�C����t�y6�@̐nՊJ�쨃L��:�P]86��Ӓ�i��YB�*�l�� ���5"L�ePc>G�']�{ɇ4D~�����w�{'�!��A�,��l���G�4������+��7;��u�AU�qK��ź*���>g������T�p�#��B%�>`R{DQ�֔
��퉰{;FJ��V7���9������m�93�ֲX�G�8�Z���������Fa��PT(L'<�f�޹��g � ��ڢ���U�90xM��١�n"�t��C'z"2oZH�]=(����W�k�;�i^(�v�dd.-nvL�p���0}<�����ނtw��hK&&��z.sJ��y�BC�Mt����l��8�J0�EB-eI:�eY��h���L:����DC*D�E�"�$�p���(�&��v-�I1��PA���%����]r{�9��;/_2�Ð����� �g�X��.ȝ%w�v�4�R͇����7�g&z�!��S��p��NEʳ�"l�sPw��Uܰ�K��B��C�eۧӮ��;|���a�(���=Y����fIwm��۵Ф�VY���p� � ��������d�B�7�<���2�͗�j���E��/��&���^�����/w�<����s"��W[�S�d^�D. �c&��c2z��V�|!��jp3M�~m��"�E��r�̩���3�5�Ҋ�GIh����>�}
;�z�yq{�(=s���|�ut�u�>���t{��i��M�m�ו5		#���@xc,��\��B�Q4 4�Y���#��_�!���� U�̒�I*L �!��X�PiU��0!���^,<�T!�jK��/!�'�� �hBcM��/c=�D�>x�2�1����̿���S���:�~�v�wS�:(Q�V8�����7�N��Rn~�~;����\�@r��9u��O�dJ��h\� P0`�$���?TR�S��lE�@�a����1wZ���1qB�
I�?c�y�3��I9Є��h��8�1 �M����A���ҽ�1�y�ř������q�=B\����3��p�F�.����@�,��	)V�-Q�ل3��ߦM�)�m^�2�������K.OXn0~��{�Pʯ��L�	0Q@�NI��8��l����N ($0'��3ŝ+�6��ܣLOIN�qL�^��\�����ɍ5�(mL� �&���a�ؔ�0uZd06�P����� �4������� ���N�9@H'�y�b<E���,9*,O mV=4�/�.H`�ƽ�M��65#$�B5TlB07�S�<�����@��*%D@��U%Z��)�!8���'�(��Rahi�P5���I&��5/�V.SP_��-�@8J�
���t�?J�<z��������V\�p�P�f6ڙ�
�*@1�r�2���Q|�H &Z�O�|6�K:��v%��H � �b���r�P�:,U*�d�)�;�Μ��M��m[�b���75��v_MF��Ψ�Hodq���˔���;���^�$Y��A�;�� UUl9T�eHA��������玌�)�[��%-v���+��b��_�G���^�堥nn�%)�����V��$]s�X0�#z�$�ͣ>��q�L�$8a1�2	V$_���"�(H&GR� 