BZh91AY&SY�sk' M߀Py���g߰����P~5څE��PR�چU4f��4h�2b� $I�h��Q�h�� P  �!$M��56��0i d�   �0L@0	�h�h`b`�$i4!��ꞣmcL�A�����h��B�I	hIxF�=�������n`xR�H��*-Q��mUh��&jCL�4*Ԗ��(�Q��q��y�G��wZ��䡍���BU8��9�^�d��J,9��eN5ٕ�{��[�]�Vz��͠���K��$.Mt����xݼ�'�/'0#%�f!
kRנ$��U:��x��Lap�|��&L�շ*Yn��J���v�6L�˅J�����^����g|�J;�$G��!�����4�+4�"�jĜ��9��$g-9�YҤMؠ�\��F�n&��=c
�kZ�y%�&���CIgTi�бSN�ӹ�Tf4a֐�06�����o�61��6�i4�!�������/�U%&���q�r�b(}�(`�ʌkKFT)��P��}�a}�E�#�(0��)��ClZZ�	�����h�Wq������^v��˘�e�y��a��^ �p�s�|��(8I��\�i$F�
0S�}E����9(N�Q?�Ȳy�T�;M�I�v��5��o�{���H�w��J�{��])�ZobZ҂�j4���m�F�����C�_�3���EȿXC�pS�+B�4�%�D0�Xm�(5��E\	e�,��TY��˟Q�u�����Ii2Ra+��6�Nm&���u#aK��ս9�3�R��ɏc���\m�����Ar�Ka�.+���[7��6,KI��M��vopi7L'�`t69[ӥȶ�����o���TW��v�������L�.V���p���N�PҮ.�WE0�n�ju�@Һ�ma�r�xŹJYf�$����D�iɂ^}���1�x���J'������./��d��-F�dzL��q����bm�^w��N�[�����|=>����8�K5$�mep:K3���`]1�vH/)�x�|(�Y$�q������JtDܞL^�}�N���sQ�F��=�=�hW�p�PT�*O�:ӀW-���+h:�+��E@��P�jXX�#Y��r�R��M��ӱ�ɚsf��V�
ҀN"�X�_�C��,�~EFkz';_{�:�����7�e)ֳ��8���9���.�p�!���N